<?xml version="1.0" encoding="utf-8"?>

<!-- - - - - - - - - - - - - - - - - - - - - - - - - - - - - -->
<!-- Electricity Networks Lib                                -->
<!--                                                         -->
<!-- This Electricity Networks Lib is made available         -->
<!-- under the Open Data Commons Attribution License:        -->
<!-- http://opendatacommons.org/licenses/by/1.0/             -->
<!--                                                         -->
<!-- If you use the data in this file please cite            -->
<!--                                                         -->
<!-- Lars Schewe, Martin Schmidt: "Electricity Networks Lib" -->
<!-- - - - - - - - - - - - - - - - - - - - - - - - - - - - - -->

<cdl>
  <info title="Grimm_et_al_2015_6_node" date="2015-11-13" author="Martin Schmidt"
	description="Network taken from the paper Grimm et al. (2015).
		     It is roughly based on the network used in Chao and Peck (1998)."/>
  <candidateLines>
    <candidateLine from="node_1" id="cand_line_1" to="node_6">
      <capacity unit="MW" value="200"/>
      <susceptance unit="S" value="0.5"/>
      <investmentCosts unit="EUR" value="230000"/>
    </candidateLine>
    <candidateLine from="node_2" id="cand_line_2" to="node_5">
      <capacity unit="MW" value="200"/>
      <susceptance unit="S" value="0.5"/>
      <investmentCosts unit="EUR" value="230000"/>
    </candidateLine>
  </candidateLines>
</cdl>
